library verilog;
use verilog.vl_types.all;
entity final_project_soc_nios2_qsys_0_nios2_performance_monitors is
end final_project_soc_nios2_qsys_0_nios2_performance_monitors;
