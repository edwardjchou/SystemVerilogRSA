library verilog;
use verilog.vl_types.all;
entity final_project_soc_mm_interconnect_0 is
    port(
        clk_0_clk_clk   : in     vl_logic;
        sdram_pll_c0_clk: in     vl_logic;
        nios2_qsys_0_reset_n_reset_bridge_in_reset_reset: in     vl_logic;
        sdram_reset_reset_bridge_in_reset_reset: in     vl_logic;
        nios2_qsys_0_data_master_address: in     vl_logic_vector(25 downto 0);
        nios2_qsys_0_data_master_waitrequest: out    vl_logic;
        nios2_qsys_0_data_master_byteenable: in     vl_logic_vector(3 downto 0);
        nios2_qsys_0_data_master_read: in     vl_logic;
        nios2_qsys_0_data_master_readdata: out    vl_logic_vector(31 downto 0);
        nios2_qsys_0_data_master_write: in     vl_logic;
        nios2_qsys_0_data_master_writedata: in     vl_logic_vector(31 downto 0);
        nios2_qsys_0_data_master_debugaccess: in     vl_logic;
        nios2_qsys_0_instruction_master_address: in     vl_logic_vector(25 downto 0);
        nios2_qsys_0_instruction_master_waitrequest: out    vl_logic;
        nios2_qsys_0_instruction_master_read: in     vl_logic;
        nios2_qsys_0_instruction_master_readdata: out    vl_logic_vector(31 downto 0);
        jtag_uart_0_avalon_jtag_slave_address: out    vl_logic_vector(0 downto 0);
        jtag_uart_0_avalon_jtag_slave_write: out    vl_logic;
        jtag_uart_0_avalon_jtag_slave_read: out    vl_logic;
        jtag_uart_0_avalon_jtag_slave_readdata: in     vl_logic_vector(31 downto 0);
        jtag_uart_0_avalon_jtag_slave_writedata: out    vl_logic_vector(31 downto 0);
        jtag_uart_0_avalon_jtag_slave_waitrequest: in     vl_logic;
        jtag_uart_0_avalon_jtag_slave_chipselect: out    vl_logic;
        led_s1_address  : out    vl_logic_vector(1 downto 0);
        led_s1_write    : out    vl_logic;
        led_s1_readdata : in     vl_logic_vector(31 downto 0);
        led_s1_writedata: out    vl_logic_vector(31 downto 0);
        led_s1_chipselect: out    vl_logic;
        nios2_qsys_0_jtag_debug_module_address: out    vl_logic_vector(8 downto 0);
        nios2_qsys_0_jtag_debug_module_write: out    vl_logic;
        nios2_qsys_0_jtag_debug_module_read: out    vl_logic;
        nios2_qsys_0_jtag_debug_module_readdata: in     vl_logic_vector(31 downto 0);
        nios2_qsys_0_jtag_debug_module_writedata: out    vl_logic_vector(31 downto 0);
        nios2_qsys_0_jtag_debug_module_byteenable: out    vl_logic_vector(3 downto 0);
        nios2_qsys_0_jtag_debug_module_waitrequest: in     vl_logic;
        nios2_qsys_0_jtag_debug_module_debugaccess: out    vl_logic;
        onchip_memory2_0_s1_address: out    vl_logic_vector(1 downto 0);
        onchip_memory2_0_s1_write: out    vl_logic;
        onchip_memory2_0_s1_readdata: in     vl_logic_vector(31 downto 0);
        onchip_memory2_0_s1_writedata: out    vl_logic_vector(31 downto 0);
        onchip_memory2_0_s1_byteenable: out    vl_logic_vector(3 downto 0);
        onchip_memory2_0_s1_chipselect: out    vl_logic;
        onchip_memory2_0_s1_clken: out    vl_logic;
        sdram_s1_address: out    vl_logic_vector(22 downto 0);
        sdram_s1_write  : out    vl_logic;
        sdram_s1_read   : out    vl_logic;
        sdram_s1_readdata: in     vl_logic_vector(15 downto 0);
        sdram_s1_writedata: out    vl_logic_vector(15 downto 0);
        sdram_s1_byteenable: out    vl_logic_vector(1 downto 0);
        sdram_s1_readdatavalid: in     vl_logic;
        sdram_s1_waitrequest: in     vl_logic;
        sdram_s1_chipselect: out    vl_logic;
        sdram_pll_pll_slave_address: out    vl_logic_vector(1 downto 0);
        sdram_pll_pll_slave_write: out    vl_logic;
        sdram_pll_pll_slave_read: out    vl_logic;
        sdram_pll_pll_slave_readdata: in     vl_logic_vector(31 downto 0);
        sdram_pll_pll_slave_writedata: out    vl_logic_vector(31 downto 0);
        sysid_qsys_0_control_slave_address: out    vl_logic_vector(0 downto 0);
        sysid_qsys_0_control_slave_readdata: in     vl_logic_vector(31 downto 0);
        to_hw_port_s1_address: out    vl_logic_vector(1 downto 0);
        to_hw_port_s1_write: out    vl_logic;
        to_hw_port_s1_readdata: in     vl_logic_vector(31 downto 0);
        to_hw_port_s1_writedata: out    vl_logic_vector(31 downto 0);
        to_hw_port_s1_chipselect: out    vl_logic;
        to_hw_sig_s1_address: out    vl_logic_vector(1 downto 0);
        to_hw_sig_s1_write: out    vl_logic;
        to_hw_sig_s1_readdata: in     vl_logic_vector(31 downto 0);
        to_hw_sig_s1_writedata: out    vl_logic_vector(31 downto 0);
        to_hw_sig_s1_chipselect: out    vl_logic;
        to_sw_port_s1_address: out    vl_logic_vector(1 downto 0);
        to_sw_port_s1_readdata: in     vl_logic_vector(31 downto 0);
        to_sw_sig_s1_address: out    vl_logic_vector(1 downto 0);
        to_sw_sig_s1_readdata: in     vl_logic_vector(31 downto 0)
    );
end final_project_soc_mm_interconnect_0;
