library verilog;
use verilog.vl_types.all;
entity testbench_gend is
end testbench_gend;
